module Not(A,O);

    input A;
    output O;

    assign O = ~A;

endmodule